library verilog;
use verilog.vl_types.all;
entity des3 is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        x               : out    vl_logic
    );
end des3;
