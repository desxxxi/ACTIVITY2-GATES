library verilog;
use verilog.vl_types.all;
entity des51_tb is
end des51_tb;
