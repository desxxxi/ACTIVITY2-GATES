library verilog;
use verilog.vl_types.all;
entity des4 is
    port(
        x               : in     vl_logic;
        y               : in     vl_logic;
        z               : in     vl_logic;
        m               : out    vl_logic
    );
end des4;
