library verilog;
use verilog.vl_types.all;
entity des3_tb is
end des3_tb;
