library verilog;
use verilog.vl_types.all;
entity des2_tb is
end des2_tb;
