library verilog;
use verilog.vl_types.all;
entity des1_tb is
end des1_tb;
