library verilog;
use verilog.vl_types.all;
entity des51 is
    port(
        d0              : in     vl_logic;
        d1              : in     vl_logic;
        s               : in     vl_logic;
        a               : out    vl_logic
    );
end des51;
