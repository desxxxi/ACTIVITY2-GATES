library verilog;
use verilog.vl_types.all;
entity des52_tb is
end des52_tb;
