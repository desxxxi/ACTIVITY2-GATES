library verilog;
use verilog.vl_types.all;
entity des1 is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        d               : in     vl_logic;
        e               : out    vl_logic
    );
end des1;
