library verilog;
use verilog.vl_types.all;
entity des2 is
    port(
        i               : in     vl_logic;
        m               : in     vl_logic;
        r               : in     vl_logic;
        l               : in     vl_logic;
        e               : out    vl_logic
    );
end des2;
