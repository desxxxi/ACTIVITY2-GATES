library verilog;
use verilog.vl_types.all;
entity des4_tb is
end des4_tb;
