library verilog;
use verilog.vl_types.all;
entity des53_tb is
end des53_tb;
